// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);

/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

    // Address decoding: Each SRAM gets 64KB (16384 words * 4 bytes = 65536 bytes)
    // SRAM 0: 0x00000000 - 0x0000FFFF
    // SRAM 1: 0x00010000 - 0x0001FFFF
    // SRAM 2: 0x00020000 - 0x0002FFFF
    wire [1:0] sram_sel;
    assign sram_sel = wbs_adr_i[17:16];  // Upper 2 bits of address select which SRAM

    // Internal signals for each SRAM instance
    wire wbs_ack_o_0, wbs_ack_o_1, wbs_ack_o_2;
    wire [31:0] wbs_dat_o_0, wbs_dat_o_1, wbs_dat_o_2;
    wire wbs_stb_i_0, wbs_stb_i_1, wbs_stb_i_2;

    // Address decoding: only assert strobe for the selected SRAM
    assign wbs_stb_i_0 = wbs_stb_i && (sram_sel == 2'b00);
    assign wbs_stb_i_1 = wbs_stb_i && (sram_sel == 2'b01);
    assign wbs_stb_i_2 = wbs_stb_i && (sram_sel == 2'b10);

    // Combine acknowledge signals
    assign wbs_ack_o = wbs_ack_o_0 | wbs_ack_o_1 | wbs_ack_o_2;

    // Multiplex data outputs based on which SRAM responded
    assign wbs_dat_o = (sram_sel == 2'b00) ? wbs_dat_o_0 :
                       (sram_sel == 2'b01) ? wbs_dat_o_1 :
                       (sram_sel == 2'b10) ? wbs_dat_o_2 : 32'b0;

    // SRAM instance 0 (base address)
    CF_SRAM_16384x32 sram (
    `ifdef USE_POWER_PINS
        .VPWR(vccd1),   // User area 1 1.8V power
        .VGND(vssd1),   // User area 1 digital ground
    `endif

        // Wishbone Bus Interface
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .wbs_stb_i(wbs_stb_i_0),
        .wbs_cyc_i(wbs_cyc_i),
        .wbs_we_i(wbs_we_i),
        .wbs_sel_i(wbs_sel_i),
        .wbs_dat_i(wbs_dat_i),
        .wbs_adr_i(wbs_adr_i[15:0]),  // Lower 16 bits for 64KB address space
        .wbs_ack_o(wbs_ack_o_0),
        .wbs_dat_o(wbs_dat_o_0)
    );

    // SRAM instance 1 (offset 0x10000)
    CF_SRAM_16384x32 sram1 (
    `ifdef USE_POWER_PINS
        .VPWR(vccd1),   // User area 1 1.8V power
        .VGND(vssd1),   // User area 1 digital ground
    `endif

        // Wishbone Bus Interface
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .wbs_stb_i(wbs_stb_i_1),
        .wbs_cyc_i(wbs_cyc_i),
        .wbs_we_i(wbs_we_i),
        .wbs_sel_i(wbs_sel_i),
        .wbs_dat_i(wbs_dat_i),
        .wbs_adr_i(wbs_adr_i[15:0]),  // Lower 16 bits for 64KB address space
        .wbs_ack_o(wbs_ack_o_1),
        .wbs_dat_o(wbs_dat_o_1)
    );

    // SRAM instance 2 (offset 0x20000)
    CF_SRAM_16384x32 sram2 (
    `ifdef USE_POWER_PINS
        .VPWR(vccd1),   // User area 1 1.8V power
        .VGND(vssd1),   // User area 1 digital ground
    `endif

        // Wishbone Bus Interface
        .wb_clk_i(wb_clk_i),
        .wb_rst_i(wb_rst_i),
        .wbs_stb_i(wbs_stb_i_2),
        .wbs_cyc_i(wbs_cyc_i),
        .wbs_we_i(wbs_we_i),
        .wbs_sel_i(wbs_sel_i),
        .wbs_dat_i(wbs_dat_i),
        .wbs_adr_i(wbs_adr_i[15:0]),  // Lower 16 bits for 64KB address space
        .wbs_ack_o(wbs_ack_o_2),
        .wbs_dat_o(wbs_dat_o_2)
    );

// Tie off unused outputs
assign la_data_out = 128'b0;
assign io_out = {`MPRJ_IO_PADS{1'b0}};
assign io_oeb = {`MPRJ_IO_PADS{1'b1}};  // Set all IOs as inputs (output enable bar = 1)
assign user_irq = 3'b0;

endmodule	// user_project_wrapper

`default_nettype wire
